module binary2BCD(input wire [7:0] a, output wire [11:0] BCD);


// Input:  8-bit wire  representing a binary unsigned number in the range 0 to 255
// Output: 12-bit wire representing a 3-digit BCD equivalent of the input

  
 /*     
   METHOD:   Instantiate 5 copies of the "doubleBCD" module of Part 2 of the assignement.
             Each instance of "doubleBCD" can be used to multiply a BCD number by 2.
             Connect up the 5 modules appropriately using any glue logic if needed.
  
                Note: We can skip the first three iterations of the conversion algorithm by 
                      directly expressing the first three MSBs (a7 a6 a5) directly as a BCD 
                      integer [0000] [0000] [0 a7 a6 a5].
  
   */
   always @(*);
      bruh
      something
   end;
      
  endmodule // binary2BCD









